`ifndef __CONTAINER_PKG_SV__
`define __CONTAINER_PKG_SV__
package container_pkg;
  `include  "base_iterator.svh"
  `include  "container.svh"
  `include  "container_utility_macros.svh"

  `include  "array.svh"
  `include  "ordered_map.svh"

  `include  "container_manipulation_macros.svh"
endpackage
`endif
